module rtfhiewfbwhejbfewbfewbfuewfl;
endmodule
