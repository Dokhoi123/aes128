module rtl;
endmodule
