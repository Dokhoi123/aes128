module sub_bytes
