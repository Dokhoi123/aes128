module sub_bytes( 
input  
